module tb1();
